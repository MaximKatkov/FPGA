	
	module IP_example_test;
 
	IP_example_tb IP_example_task();
  
		initial
			begin
		    
				IP_example_task.reset;
			
			//fork
			
			//state_machine_task.reset;
			//state_machine_task.reset;
			//state_machine_task.reset;
			//state_machine_task.reset;
			
			//join
			
			
			end

	endmodule // IP_example_task