	
	module FIFO_example_test;
 
	FIFO_example_tb FIFO_example_task();
  
		initial
			begin
		    
				FIFO_example_task.reset;
			
			end

	endmodule // FIFO_example_task