
	module CDC_test;
 
	CDC_tb CDC_task();
  
		initial
			begin
		    
				CDC_task.reset;
			
			end

	endmodule // CDC_task