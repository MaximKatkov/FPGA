
 module state_machine_test;
 
 state_machine_tb state_machine_task();
  
    initial
	    begin
		    
			state_machine_task.reset;
			
			//fork
			
			//state_machine_task.reset;
			//state_machine_task.reset;
			//state_machine_task.reset;
			//state_machine_task.reset;
			
			//join
			
			
		end

 endmodule // state_machine_task