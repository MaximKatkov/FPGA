/**************************************************************************************************  
 *                                                                                                *
 *  File Name:     rkob_ptp_ram.v         		        									      *
 *                                                                                                *
 **************************************************************************************************
 *                                                                                                *
 *  Description:   Version P2P                 				                                      *
 *                                                                                                *
 *                                                                                                *
 *                                                                                                *
 **************************************************************************************************
 *  Verilog Code                                                                                  *
 **************************************************************************************************/
 
 module rkob_ptp_ram (clk, we, wr_addr, rd_addr, wr_data, rd_data);

/**************************************************************************************************
 *      PARAMETERS                                                                                *
 **************************************************************************************************/
 
 parameter DATA_WIDTH = 52; 
 parameter ADDR_WIDTH = 12; 
 parameter MEM_DEPTH  = 4096;
 
/**************************************************************************************************
 *      INPUT PORTS                                                                               *
 **************************************************************************************************/ 
 
 input 						clk;
 input 						we;
 
 input 	[ADDR_WIDTH - 1:0] 	wr_addr;
 input 	[ADDR_WIDTH - 1:0] 	rd_addr;
 
 input  [DATA_WIDTH - 1:0] 	wr_data;
 
/**************************************************************************************************
 *      OUTPUT PORTS                                                                              *
 **************************************************************************************************/
  
 output [DATA_WIDTH - 1:0] 	rd_data;

/**************************************************************************************************
 *      WIRES & REGS                                                                              *
 **************************************************************************************************/ 
 
 reg 	[DATA_WIDTH - 1:0] 	ram [MEM_DEPTH - 1:0];
 reg 	[ADDR_WIDTH - 1:0] 	rd_addr_r;

/**************************************************************************************************
 *      CONTENT                                                                                   *
 **************************************************************************************************/ 
 
 integer i;                                        // Обнулим все ячейки памяти
 initial
	begin
		for (i = 0; i < MEM_DEPTH; i = i + 1)
			begin
				ram[i] = {(DATA_WIDTH){1'b0}};					
			end	
	end

 always @(posedge clk) 
    begin
        if (we)
            ram[wr_addr] <= wr_data;
      
         rd_addr_r <= rd_addr;
     end
     
 assign rd_data = ram[rd_addr_r];

 endmodule // rkob_ptp_ram
